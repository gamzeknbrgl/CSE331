`define DELAY 20
module mux_2x1_32_bit_testbench();
reg[31:0]d0;
reg[31:0]d1;
reg s;

wire [31:0]outp;

mux_2x1_32_bit result(outp,d0,d1,s);

initial begin
d0=32'b00000000000000000000000000000011; d1=32'b00000000000000000000000000000001; s=1'b1;
#`DELAY;
d0=32'b00000000000000000000000000000010; d1=32'b0100000000000000000000000000001; s=1'b0;
#`DELAY;
d0=32'b11111111111111111111111111111111; d1=32'b11111111111111111111111111111111; s=1'b0;
#`DELAY;
d0=32'b01111111111111111111111111111111; d1=32'b0000000000000000000000000000001; s=1'b1;
#`DELAY;
d0=32'b00000000000000000000000000111111; d1=32'b0000000000000000000000000111011; s=1'b0;
end
initial begin
$monitor("time=%2d, d0=%32b, d1=%32b, s=%1b, output=%32b",$time,d0,d1,s,outp);
end

endmodule