`define DELAY 20
module full_adder_32_bit_testbench();
reg [31:0]a,b;
reg c_in;
wire [31:0]sum;
wire c_out;
full_adder_32_bit fa32b(sum,c_out,a,b,c_in);

initial begin
a=32'b00000000000000000000000000000011; b=32'b00000000000000000000000000000001; c_in=1'b1;
#`DELAY;
a=32'b00000000000000000000000000000010; b=32'b0100000000000000000000000000001; c_in=1'b0;
#`DELAY;
a=32'b11111111111111111111111111111111; b=32'b11111111111111111111111111111111; c_in=1'b0;
#`DELAY;
a=32'b01111111111111111111111111111111; b=32'b0000000000000000000000000000001; c_in=1'b0;
#`DELAY;
a=32'b00000000000000000000000000111111; b=32'b0000000000000000000000000111111; c_in=1'b0;
end
initial begin
$monitor("time=%2d, a=%32b, b=%32b, c_in=%1b, sum=%32b, c_out=%1b",$time,a,b,c_in,sum,c_out);
end

endmodule