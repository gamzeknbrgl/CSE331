`define DELAY 20
module myXor_32bit_testbench();
reg [31:0]a,b;
wire [31:0]out;

myXor_32bit xor_32bit(out,a,b);

initial begin
a=32'b00000000000000000000000000000011; b=32'b00000000000000000000000000000001; 
#`DELAY;
a=32'b00000000000000000000000000000010; b=32'b0100000000000000000000000000001; 
#`DELAY;
a=32'b11111111111111111111111111111111; b=32'b11111111111111111111111111111111; 
#`DELAY;
a=32'b01111111111111111111111111111111; b=32'b0000000000000000000000000000001; 
#`DELAY;
a=32'b00000000000000000000000000111111; b=32'b0000000000000000000000000111111; 
end
initial begin
$monitor("time=%2d, a=%32b, b=%32b, output=%32b",$time,a,b,out);
end

endmodule