`define DELAY 20
module ALU_32Bit_testbench(); 
reg [31:0]ai;
reg [31:0]bi;
reg aluop0, aluop1, aluop2,  cin;
wire [31:0]outp;
wire cout;

ALU_32Bit a1(outp,cout, aluop0, aluop1, aluop2, ai,bi, cin);

initial begin
$display("Test Results");
$display("And:");
ai = 32'b00000000000000000000000000000000; bi = 32'b00000000000000000000000000000000; aluop0= 1'b0; aluop1= 1'b0; aluop2= 1'b0; cin= 1'b0; 
#`DELAY;
ai = 32'b00000000000000000000000000000001; bi = 32'b00000000000000000000000000000000; aluop0= 1'b0; aluop1= 1'b0; aluop2= 1'b0; cin= 1'b0;
#`DELAY;
ai = 32'b00000000000000000000000000000000; bi = 32'b00000000000000000000000000000001; aluop0= 1'b0; aluop1= 1'b0; aluop2= 1'b0; cin= 1'b0;  
#`DELAY;
ai = 32'b11111111111111111111111111111111; bi = 32'b11111111111111111111111111111111; aluop0= 1'b0; aluop1= 1'b0; aluop2= 1'b0; cin= 1'b0;
#`DELAY;
$display("Or:");
#`DELAY;
ai = 32'b00000000000000000000000000000000; bi = 32'b00000000000000000000000000000000; aluop0= 1'b1; aluop1= 1'b0; aluop2= 1'b0; cin= 1'b0; 
#`DELAY;
ai = 32'b00000000000000000000000000000001; bi = 32'b00000000000000000000000000000000; aluop0= 1'b1; aluop1= 1'b0; aluop2= 1'b0; cin= 1'b0;
#`DELAY;
ai = 32'b00000000000000000000000000000000; bi = 32'b00000000000000000000000000000001; aluop0= 1'b1; aluop1= 1'b0; aluop2= 1'b0; cin= 1'b0;  
#`DELAY;
ai = 32'b11111111111111111111111111111111; bi = 32'b11111111111111111111111111111111; aluop0= 1'b1; aluop1= 1'b0; aluop2= 1'b0; cin= 1'b0;
#`DELAY;
$display("Add:");
#`DELAY;
ai = 32'b00000000000000000000000000000000; bi = 32'b00000000000000000000000000000000; aluop0= 1'b0; aluop1= 1'b1; aluop2= 1'b0; cin= 1'b0; 
#`DELAY;
ai = 32'b00000000000000000000000000000001; bi = 32'b00000000000000000000000000000000; aluop0= 1'b0; aluop1= 1'b1; aluop2= 1'b0; cin= 1'b0;
#`DELAY;
ai = 32'b00000000000000000000000000000000; bi = 32'b00000000000000000000000000000001; aluop0= 1'b0; aluop1= 1'b1; aluop2= 1'b0; cin= 1'b0;  
#`DELAY;
ai = 32'b11111111111111111111111111111111; bi = 32'b11111111111111111111111111111111; aluop0= 1'b0; aluop1= 1'b1; aluop2= 1'b0; cin= 1'b0;
#`DELAY;
$display("Substract:");
#`DELAY;
ai = 32'b00000000000000000000000000000000; bi = 32'b00000000000000000000000000000000; aluop0= 1'b0; aluop1= 1'b1; aluop2= 1'b1; cin= 1'b1; 
#`DELAY;
ai = 32'b00000000000000000000000000000001; bi = 32'b00000000000000000000000000000000; aluop0= 1'b0; aluop1= 1'b1; aluop2= 1'b1; cin= 1'b1;
#`DELAY;
ai = 32'b00000000000000000000000000000000; bi = 32'b00000000000000000000000000000001; aluop0= 1'b0; aluop1= 1'b1; aluop2= 1'b1; cin= 1'b1;  
#`DELAY;
ai = 32'b11111111111111111111111111111111; bi = 32'b11111111111111111111111111111111; aluop0= 1'b0; aluop1= 1'b1; aluop2= 1'b1; cin= 1'b1;
#`DELAY;
$display("Set-on-less-than:");
#`DELAY;
ai = 32'b00000000000000000000000000000000; bi = 32'b00000000000000000000000000000000; aluop0= 1'b1; aluop1= 1'b1; aluop2= 1'b1; cin= 1'b1; 
#`DELAY;
ai = 32'b00000000000000000000000000000001; bi = 32'b00000000000000000000000000000000; aluop0= 1'b1; aluop1= 1'b1; aluop2= 1'b1; cin= 1'b1;
#`DELAY;
ai = 32'b00000000000000000000000000000000; bi = 32'b00000000000000000000000000000001; aluop0= 1'b1; aluop1= 1'b1; aluop2= 1'b1; cin= 1'b1;  
#`DELAY;
ai = 32'b11111111111111111111111111111111; bi = 32'b11111111111111111111111111111111; aluop0= 1'b1; aluop1= 1'b1; aluop2= 1'b1; cin= 1'b1;
end


initial
begin
$monitor("time = %2d, ai =%32b, bi=%32b, outp=%32b, cout=%1b, cin: %1b", $time, ai, bi, outp, cout,cin );
end

 

endmodule